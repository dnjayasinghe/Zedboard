----------------------------------------------------------------------------------
--
-- Copyright 2019 Ruhr University Bochum, Horst Görtz Institute for IT Security
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy of this software
-- and associated documentation files (the "Software"), to deal in the Software without restriction, 
-- including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, 
-- and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do 
-- so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in all copies or substantial 
-- portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT 
-- LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. 
-- IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, 
-- WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE 
-- SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

------------------------------------------------------------------
-- Entity 
------------------------------------------------------------------ 
entity sbox is
	port(
		encrypt	: in std_logic;
		input		: in std_logic_vector(31 downto 0);
		output	: out std_logic_vector(31 downto 0)
		);
end entity sbox;

------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------ 
architecture dfl of sbox is

------------------------------------------------------------------
-- Components
------------------------------------------------------------------ 
component sbox8 is
	port(
		encrypt	: in std_logic;
		input		: in std_logic_vector(7 downto 0);
		output	: out std_logic_vector(7 downto 0)
		);
end component sbox8;

------------------------------------------------------------------
-- Begin
------------------------------------------------------------------ 
begin

	bits31_24: sbox8
	port map(
		encrypt => encrypt,
		input => input(31 downto 24),
		output => output(31 downto 24));
		
	bits23_16: sbox8
	port map(
		encrypt => encrypt,
		input => input(23 downto 16),
		output => output(23 downto 16));
		
	bits15_8: sbox8
	port map(
		encrypt => encrypt,
		input => input(15 downto 8),
		output => output(15 downto 8));
		
	bits7_0: sbox8
	port map(
		encrypt => encrypt,
		input => input(7 downto 0),
		output => output(7 downto 0));

end architecture;